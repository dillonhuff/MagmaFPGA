

module top(
	input [0 : 0] in_wire_0,
	input [0 : 0] in_wire_1,
	input [31 : 0] config_addr,
	input [0 : 0] clk,
	input [0 : 0] in_wire_2,
	input [0 : 0] reset,
	input [31 : 0] config_data,
	output [0 : 0] out_wire_0,
	output [0 : 0] out_wire_1,
	output [0 : 0] out_wire_2
	);

	// Internal wires
/* verilator lint_off PINMISSING */

	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_18;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_36;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_0_1_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_side_1_track_3_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_1_pin_1_to_pe_tile_2_1_side_1_track_1_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_side_1_track_1_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_0side_2_track_0_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_0;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] out_pad_1_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_26;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_0_pin_1_to_pe_tile_2_0_side_1_track_1_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_10;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_1_0_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_0_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_0side_2_track_3_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0_side_1_track_2_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_1_pin_3_to_pe_tile_2_1_side_1_track_3_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_32;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_2_pin_1_to_pe_tile_0_2_side_3_track_1_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_0_pin_0_to_pe_tile_0_0_side_3_track_0_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_43;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_21;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_35;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_2_2_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_25;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_1_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_41;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_2_const;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_42;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_47;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0_side_1_track_1_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_1_pin_2_to_pe_tile_0_1_side_3_track_2_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0side_2_track_0_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_1;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_33;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_0_pin_3_to_pe_tile_2_0_side_1_track_3_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_2_pin_3_to_pe_tile_2_2_side_1_track_3_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_16;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_3_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_1_side_1_track_1_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_0_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_1_side_1_track_2_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_9;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_2_pin_1_to_pe_tile_2_2_side_1_track_1_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_0side_2_track_0_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_1_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_28;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_2_pin_2_to_pe_tile_2_2_side_1_track_2_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_11;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_46;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_1_pin_1_to_pe_tile_0_1_side_3_track_1_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_6;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_3;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_19;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_38;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_13;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_2;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_0_0_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_0_pin_1_to_pe_tile_0_0_side_3_track_1_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_5;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_7;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_15;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_3;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_2_0_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_2_1_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_31;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_4;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0side_2_track_3_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_45;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_2_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_1_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_0side_2_track_2_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_0side_2_track_3_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_side_1_track_2_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_2_pin_3_to_pe_tile_0_2_side_3_track_3_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_1_pin_0_to_pe_tile_2_1_side_1_track_0_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_34;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_side_1_track_0_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_1_side_1_track_0_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_24;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_0_pin_2_to_pe_tile_0_0_side_3_track_2_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_27;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_29;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_0side_2_track_1_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_0_pin_2_to_pe_tile_2_0_side_1_track_2_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0_side_1_track_0_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_1_side_1_track_3_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_14;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_0_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_20;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_3;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_0_2_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_1_2_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_30;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_2_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_12;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_0_pin_3_to_pe_tile_0_0_side_3_track_3_in;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] out_pad_0_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] wire_8;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_3_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0_side_1_track_3_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0side_2_track_1_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_0_pin_0_to_pe_tile_2_0_side_1_track_0_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_40;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_37;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_22;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_23;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_1_pin_3_to_pe_tile_0_1_side_3_track_3_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_2_pin_0_to_pe_tile_2_2_side_1_track_0_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_44;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_2_0side_2_track_2_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_2_pin_2_to_pe_tile_0_2_side_3_track_2_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_2_pin_0_to_pe_tile_0_2_side_3_track_0_in;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_39;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] wire_17;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_1;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_2;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_0_0side_2_track_1_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] in_pad_1_pin_0_to_pe_tile_0_1_side_3_track_0_in;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] out_pad_2_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_3_const;
	/* verilator lint_off UNOPTFLAT */
	wire [16 - 1 : 0] pe_tile_1_1_id_wire;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_3;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] pe_tile_1_0side_2_track_2_in_const;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] out_pad_1_pin_2_to_pe_tile_2_1_side_1_track_2_out;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_0;
	/* verilator lint_off UNOPTFLAT */
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_2;
	// End of wire declarations

	io1in_pad in_pad_0(
		.clk(clk),
		.top_pin(in_wire_0),
		.pin_0(in_pad_0_pin_0_to_pe_tile_0_0_side_3_track_0_in),
		.pin_1(in_pad_0_pin_1_to_pe_tile_0_0_side_3_track_1_in),
		.pin_2(in_pad_0_pin_2_to_pe_tile_0_0_side_3_track_2_in),
		.pin_3(in_pad_0_pin_3_to_pe_tile_0_0_side_3_track_3_in)
	);

	io1in_pad in_pad_1(
		.clk(clk),
		.top_pin(in_wire_1),
		.pin_0(in_pad_1_pin_0_to_pe_tile_0_1_side_3_track_0_in),
		.pin_1(in_pad_1_pin_1_to_pe_tile_0_1_side_3_track_1_in),
		.pin_2(in_pad_1_pin_2_to_pe_tile_0_1_side_3_track_2_in),
		.pin_3(in_pad_1_pin_3_to_pe_tile_0_1_side_3_track_3_in)
	);

	io1in_pad in_pad_2(
		.clk(clk),
		.top_pin(in_wire_2),
		.pin_0(in_pad_2_pin_0_to_pe_tile_0_2_side_3_track_0_in),
		.pin_1(in_pad_2_pin_1_to_pe_tile_0_2_side_3_track_1_in),
		.pin_2(in_pad_2_pin_2_to_pe_tile_0_2_side_3_track_2_in),
		.pin_3(in_pad_2_pin_3_to_pe_tile_0_2_side_3_track_3_in)
	);

	io1out_pad out_pad_0(
		.top_pin(out_wire_0),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(out_pad_0_id_wire),
		.pin_0(out_pad_0_pin_0_to_pe_tile_2_0_side_1_track_0_out),
		.pin_1(out_pad_0_pin_1_to_pe_tile_2_0_side_1_track_1_out),
		.pin_2(out_pad_0_pin_2_to_pe_tile_2_0_side_1_track_2_out),
		.pin_3(out_pad_0_pin_3_to_pe_tile_2_0_side_1_track_3_out)
	);

	assign_mod #(.width(16))  assign_out_pad_0_id_wire_0(
		.out(out_pad_0_id_wire),
		.in(wire_0)
	);

	const_mod #(.value(1), .width(16))  assign_out_pad_0_id_wire_0_const(
		.out(wire_0)
	);

	io1out_pad out_pad_1(
		.top_pin(out_wire_1),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(out_pad_1_id_wire),
		.pin_0(out_pad_1_pin_0_to_pe_tile_2_1_side_1_track_0_out),
		.pin_1(out_pad_1_pin_1_to_pe_tile_2_1_side_1_track_1_out),
		.pin_2(out_pad_1_pin_2_to_pe_tile_2_1_side_1_track_2_out),
		.pin_3(out_pad_1_pin_3_to_pe_tile_2_1_side_1_track_3_out)
	);

	assign_mod #(.width(16))  assign_out_pad_1_id_wire_1(
		.out(out_pad_1_id_wire),
		.in(wire_1)
	);

	const_mod #(.value(2), .width(16))  assign_out_pad_1_id_wire_1_const(
		.out(wire_1)
	);

	io1out_pad out_pad_2(
		.top_pin(out_wire_2),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(out_pad_2_id_wire),
		.pin_0(out_pad_2_pin_0_to_pe_tile_2_2_side_1_track_0_out),
		.pin_1(out_pad_2_pin_1_to_pe_tile_2_2_side_1_track_1_out),
		.pin_2(out_pad_2_pin_2_to_pe_tile_2_2_side_1_track_2_out),
		.pin_3(out_pad_2_pin_3_to_pe_tile_2_2_side_1_track_3_out)
	);

	assign_mod #(.width(16))  assign_out_pad_2_id_wire_2(
		.out(out_pad_2_id_wire),
		.in(wire_2)
	);

	const_mod #(.value(3), .width(16))  assign_out_pad_2_id_wire_2_const(
		.out(wire_2)
	);

	pe_tile pe_tile_0_0(
		.side_3_track_0_in(in_pad_0_pin_0_to_pe_tile_0_0_side_3_track_0_in),
		.side_3_track_1_in(in_pad_0_pin_1_to_pe_tile_0_0_side_3_track_1_in),
		.side_3_track_2_in(in_pad_0_pin_2_to_pe_tile_0_0_side_3_track_2_in),
		.side_3_track_3_in(in_pad_0_pin_3_to_pe_tile_0_0_side_3_track_3_in),
		.side_1_track_0_out(vertical_tile_0_0_to_tile_1_0_0),
		.side_1_track_1_out(vertical_tile_0_0_to_tile_1_0_1),
		.side_1_track_2_out(vertical_tile_0_0_to_tile_1_0_2),
		.side_1_track_3_out(vertical_tile_0_0_to_tile_1_0_3),
		.side_1_track_0_in(vertical_tile_1_0_to_tile_0_0_0),
		.side_1_track_1_in(vertical_tile_1_0_to_tile_0_0_1),
		.side_1_track_2_in(vertical_tile_1_0_to_tile_0_0_2),
		.side_1_track_3_in(vertical_tile_1_0_to_tile_0_0_3),
		.side_2_track_0_in(pe_tile_0_0side_2_track_0_in_const),
		.side_2_track_1_in(pe_tile_0_0side_2_track_1_in_const),
		.side_2_track_2_in(pe_tile_0_0side_2_track_2_in_const),
		.side_2_track_3_in(pe_tile_0_0side_2_track_3_in_const),
		.side_0_track_0_out(horizontal_tile_0_0_to_tile_0_1_0),
		.side_0_track_1_out(horizontal_tile_0_0_to_tile_0_1_1),
		.side_0_track_2_out(horizontal_tile_0_0_to_tile_0_1_2),
		.side_0_track_3_out(horizontal_tile_0_0_to_tile_0_1_3),
		.side_0_track_0_in(horizontal_tile_0_1_to_tile_0_0_0),
		.side_0_track_1_in(horizontal_tile_0_1_to_tile_0_0_1),
		.side_0_track_2_in(horizontal_tile_0_1_to_tile_0_0_2),
		.side_0_track_3_in(horizontal_tile_0_1_to_tile_0_0_3),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_0_0_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0side_2_track_0_in_const_3(
		.out(pe_tile_0_0side_2_track_0_in_const),
		.in(wire_3)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_0side_2_track_0_in_const_3_const(
		.out(wire_3)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0side_2_track_1_in_const_4(
		.out(pe_tile_0_0side_2_track_1_in_const),
		.in(wire_4)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_0side_2_track_1_in_const_4_const(
		.out(wire_4)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0side_2_track_2_in_const_5(
		.out(pe_tile_0_0side_2_track_2_in_const),
		.in(wire_5)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_0side_2_track_2_in_const_5_const(
		.out(wire_5)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0side_2_track_3_in_const_6(
		.out(pe_tile_0_0side_2_track_3_in_const),
		.in(wire_6)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_0side_2_track_3_in_const_6_const(
		.out(wire_6)
	);

	assign_mod #(.width(16))  assign_pe_tile_0_0_id_wire_7(
		.out(pe_tile_0_0_id_wire),
		.in(wire_7)
	);

	const_mod #(.value(16'd4), .width(16))  assign_pe_tile_0_0_id_wire_7_const(
		.out(wire_7)
	);

	pe_tile pe_tile_0_1(
		.side_3_track_0_in(in_pad_1_pin_0_to_pe_tile_0_1_side_3_track_0_in),
		.side_3_track_1_in(in_pad_1_pin_1_to_pe_tile_0_1_side_3_track_1_in),
		.side_3_track_2_in(in_pad_1_pin_2_to_pe_tile_0_1_side_3_track_2_in),
		.side_3_track_3_in(in_pad_1_pin_3_to_pe_tile_0_1_side_3_track_3_in),
		.side_1_track_0_out(vertical_tile_0_1_to_tile_1_1_0),
		.side_1_track_1_out(vertical_tile_0_1_to_tile_1_1_1),
		.side_1_track_2_out(vertical_tile_0_1_to_tile_1_1_2),
		.side_1_track_3_out(vertical_tile_0_1_to_tile_1_1_3),
		.side_1_track_0_in(vertical_tile_1_1_to_tile_0_1_0),
		.side_1_track_1_in(vertical_tile_1_1_to_tile_0_1_1),
		.side_1_track_2_in(vertical_tile_1_1_to_tile_0_1_2),
		.side_1_track_3_in(vertical_tile_1_1_to_tile_0_1_3),
		.side_2_track_0_out(horizontal_tile_0_1_to_tile_0_0_0),
		.side_2_track_1_out(horizontal_tile_0_1_to_tile_0_0_1),
		.side_2_track_2_out(horizontal_tile_0_1_to_tile_0_0_2),
		.side_2_track_3_out(horizontal_tile_0_1_to_tile_0_0_3),
		.side_2_track_0_in(horizontal_tile_0_0_to_tile_0_1_0),
		.side_2_track_1_in(horizontal_tile_0_0_to_tile_0_1_1),
		.side_2_track_2_in(horizontal_tile_0_0_to_tile_0_1_2),
		.side_2_track_3_in(horizontal_tile_0_0_to_tile_0_1_3),
		.side_0_track_0_out(horizontal_tile_0_1_to_tile_0_2_0),
		.side_0_track_1_out(horizontal_tile_0_1_to_tile_0_2_1),
		.side_0_track_2_out(horizontal_tile_0_1_to_tile_0_2_2),
		.side_0_track_3_out(horizontal_tile_0_1_to_tile_0_2_3),
		.side_0_track_0_in(horizontal_tile_0_2_to_tile_0_1_0),
		.side_0_track_1_in(horizontal_tile_0_2_to_tile_0_1_1),
		.side_0_track_2_in(horizontal_tile_0_2_to_tile_0_1_2),
		.side_0_track_3_in(horizontal_tile_0_2_to_tile_0_1_3),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_0_1_id_wire)
	);

	assign_mod #(.width(16))  assign_pe_tile_0_1_id_wire_8(
		.out(pe_tile_0_1_id_wire),
		.in(wire_8)
	);

	const_mod #(.value(16'd5), .width(16))  assign_pe_tile_0_1_id_wire_8_const(
		.out(wire_8)
	);

	pe_tile pe_tile_0_2(
		.side_3_track_0_in(in_pad_2_pin_0_to_pe_tile_0_2_side_3_track_0_in),
		.side_3_track_1_in(in_pad_2_pin_1_to_pe_tile_0_2_side_3_track_1_in),
		.side_3_track_2_in(in_pad_2_pin_2_to_pe_tile_0_2_side_3_track_2_in),
		.side_3_track_3_in(in_pad_2_pin_3_to_pe_tile_0_2_side_3_track_3_in),
		.side_1_track_0_out(vertical_tile_0_2_to_tile_1_2_0),
		.side_1_track_1_out(vertical_tile_0_2_to_tile_1_2_1),
		.side_1_track_2_out(vertical_tile_0_2_to_tile_1_2_2),
		.side_1_track_3_out(vertical_tile_0_2_to_tile_1_2_3),
		.side_1_track_0_in(vertical_tile_1_2_to_tile_0_2_0),
		.side_1_track_1_in(vertical_tile_1_2_to_tile_0_2_1),
		.side_1_track_2_in(vertical_tile_1_2_to_tile_0_2_2),
		.side_1_track_3_in(vertical_tile_1_2_to_tile_0_2_3),
		.side_2_track_0_out(horizontal_tile_0_2_to_tile_0_1_0),
		.side_2_track_1_out(horizontal_tile_0_2_to_tile_0_1_1),
		.side_2_track_2_out(horizontal_tile_0_2_to_tile_0_1_2),
		.side_2_track_3_out(horizontal_tile_0_2_to_tile_0_1_3),
		.side_2_track_0_in(horizontal_tile_0_1_to_tile_0_2_0),
		.side_2_track_1_in(horizontal_tile_0_1_to_tile_0_2_1),
		.side_2_track_2_in(horizontal_tile_0_1_to_tile_0_2_2),
		.side_2_track_3_in(horizontal_tile_0_1_to_tile_0_2_3),
		.side_0_track_0_in(pe_tile_0_2_in_wire_0_0_const),
		.side_0_track_1_in(pe_tile_0_2_in_wire_0_1_const),
		.side_0_track_2_in(pe_tile_0_2_in_wire_0_2_const),
		.side_0_track_3_in(pe_tile_0_2_in_wire_0_3_const),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_0_2_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_0_const_9(
		.out(pe_tile_0_2_in_wire_0_0_const),
		.in(wire_9)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_2_in_wire_0_0_const_9_const(
		.out(wire_9)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_1_const_10(
		.out(pe_tile_0_2_in_wire_0_1_const),
		.in(wire_10)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_2_in_wire_0_1_const_10_const(
		.out(wire_10)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_2_const_11(
		.out(pe_tile_0_2_in_wire_0_2_const),
		.in(wire_11)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_2_in_wire_0_2_const_11_const(
		.out(wire_11)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_3_const_12(
		.out(pe_tile_0_2_in_wire_0_3_const),
		.in(wire_12)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_0_2_in_wire_0_3_const_12_const(
		.out(wire_12)
	);

	assign_mod #(.width(16))  assign_pe_tile_0_2_id_wire_13(
		.out(pe_tile_0_2_id_wire),
		.in(wire_13)
	);

	const_mod #(.value(16'd6), .width(16))  assign_pe_tile_0_2_id_wire_13_const(
		.out(wire_13)
	);

	pe_tile pe_tile_1_0(
		.side_3_track_0_out(vertical_tile_1_0_to_tile_0_0_0),
		.side_3_track_1_out(vertical_tile_1_0_to_tile_0_0_1),
		.side_3_track_2_out(vertical_tile_1_0_to_tile_0_0_2),
		.side_3_track_3_out(vertical_tile_1_0_to_tile_0_0_3),
		.side_3_track_0_in(vertical_tile_0_0_to_tile_1_0_0),
		.side_3_track_1_in(vertical_tile_0_0_to_tile_1_0_1),
		.side_3_track_2_in(vertical_tile_0_0_to_tile_1_0_2),
		.side_3_track_3_in(vertical_tile_0_0_to_tile_1_0_3),
		.side_1_track_0_out(vertical_tile_1_0_to_tile_2_0_0),
		.side_1_track_1_out(vertical_tile_1_0_to_tile_2_0_1),
		.side_1_track_2_out(vertical_tile_1_0_to_tile_2_0_2),
		.side_1_track_3_out(vertical_tile_1_0_to_tile_2_0_3),
		.side_1_track_0_in(vertical_tile_2_0_to_tile_1_0_0),
		.side_1_track_1_in(vertical_tile_2_0_to_tile_1_0_1),
		.side_1_track_2_in(vertical_tile_2_0_to_tile_1_0_2),
		.side_1_track_3_in(vertical_tile_2_0_to_tile_1_0_3),
		.side_2_track_0_in(pe_tile_1_0side_2_track_0_in_const),
		.side_2_track_1_in(pe_tile_1_0side_2_track_1_in_const),
		.side_2_track_2_in(pe_tile_1_0side_2_track_2_in_const),
		.side_2_track_3_in(pe_tile_1_0side_2_track_3_in_const),
		.side_0_track_0_out(horizontal_tile_1_0_to_tile_1_1_0),
		.side_0_track_1_out(horizontal_tile_1_0_to_tile_1_1_1),
		.side_0_track_2_out(horizontal_tile_1_0_to_tile_1_1_2),
		.side_0_track_3_out(horizontal_tile_1_0_to_tile_1_1_3),
		.side_0_track_0_in(horizontal_tile_1_1_to_tile_1_0_0),
		.side_0_track_1_in(horizontal_tile_1_1_to_tile_1_0_1),
		.side_0_track_2_in(horizontal_tile_1_1_to_tile_1_0_2),
		.side_0_track_3_in(horizontal_tile_1_1_to_tile_1_0_3),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_1_0_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0side_2_track_0_in_const_14(
		.out(pe_tile_1_0side_2_track_0_in_const),
		.in(wire_14)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_0side_2_track_0_in_const_14_const(
		.out(wire_14)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0side_2_track_1_in_const_15(
		.out(pe_tile_1_0side_2_track_1_in_const),
		.in(wire_15)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_0side_2_track_1_in_const_15_const(
		.out(wire_15)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0side_2_track_2_in_const_16(
		.out(pe_tile_1_0side_2_track_2_in_const),
		.in(wire_16)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_0side_2_track_2_in_const_16_const(
		.out(wire_16)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0side_2_track_3_in_const_17(
		.out(pe_tile_1_0side_2_track_3_in_const),
		.in(wire_17)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_0side_2_track_3_in_const_17_const(
		.out(wire_17)
	);

	assign_mod #(.width(16))  assign_pe_tile_1_0_id_wire_18(
		.out(pe_tile_1_0_id_wire),
		.in(wire_18)
	);

	const_mod #(.value(16'd7), .width(16))  assign_pe_tile_1_0_id_wire_18_const(
		.out(wire_18)
	);

	pe_tile pe_tile_1_1(
		.side_3_track_0_out(vertical_tile_1_1_to_tile_0_1_0),
		.side_3_track_1_out(vertical_tile_1_1_to_tile_0_1_1),
		.side_3_track_2_out(vertical_tile_1_1_to_tile_0_1_2),
		.side_3_track_3_out(vertical_tile_1_1_to_tile_0_1_3),
		.side_3_track_0_in(vertical_tile_0_1_to_tile_1_1_0),
		.side_3_track_1_in(vertical_tile_0_1_to_tile_1_1_1),
		.side_3_track_2_in(vertical_tile_0_1_to_tile_1_1_2),
		.side_3_track_3_in(vertical_tile_0_1_to_tile_1_1_3),
		.side_1_track_0_out(vertical_tile_1_1_to_tile_2_1_0),
		.side_1_track_1_out(vertical_tile_1_1_to_tile_2_1_1),
		.side_1_track_2_out(vertical_tile_1_1_to_tile_2_1_2),
		.side_1_track_3_out(vertical_tile_1_1_to_tile_2_1_3),
		.side_1_track_0_in(vertical_tile_2_1_to_tile_1_1_0),
		.side_1_track_1_in(vertical_tile_2_1_to_tile_1_1_1),
		.side_1_track_2_in(vertical_tile_2_1_to_tile_1_1_2),
		.side_1_track_3_in(vertical_tile_2_1_to_tile_1_1_3),
		.side_2_track_0_out(horizontal_tile_1_1_to_tile_1_0_0),
		.side_2_track_1_out(horizontal_tile_1_1_to_tile_1_0_1),
		.side_2_track_2_out(horizontal_tile_1_1_to_tile_1_0_2),
		.side_2_track_3_out(horizontal_tile_1_1_to_tile_1_0_3),
		.side_2_track_0_in(horizontal_tile_1_0_to_tile_1_1_0),
		.side_2_track_1_in(horizontal_tile_1_0_to_tile_1_1_1),
		.side_2_track_2_in(horizontal_tile_1_0_to_tile_1_1_2),
		.side_2_track_3_in(horizontal_tile_1_0_to_tile_1_1_3),
		.side_0_track_0_out(horizontal_tile_1_1_to_tile_1_2_0),
		.side_0_track_1_out(horizontal_tile_1_1_to_tile_1_2_1),
		.side_0_track_2_out(horizontal_tile_1_1_to_tile_1_2_2),
		.side_0_track_3_out(horizontal_tile_1_1_to_tile_1_2_3),
		.side_0_track_0_in(horizontal_tile_1_2_to_tile_1_1_0),
		.side_0_track_1_in(horizontal_tile_1_2_to_tile_1_1_1),
		.side_0_track_2_in(horizontal_tile_1_2_to_tile_1_1_2),
		.side_0_track_3_in(horizontal_tile_1_2_to_tile_1_1_3),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_1_1_id_wire)
	);

	assign_mod #(.width(16))  assign_pe_tile_1_1_id_wire_19(
		.out(pe_tile_1_1_id_wire),
		.in(wire_19)
	);

	const_mod #(.value(16'd8), .width(16))  assign_pe_tile_1_1_id_wire_19_const(
		.out(wire_19)
	);

	pe_tile pe_tile_1_2(
		.side_3_track_0_out(vertical_tile_1_2_to_tile_0_2_0),
		.side_3_track_1_out(vertical_tile_1_2_to_tile_0_2_1),
		.side_3_track_2_out(vertical_tile_1_2_to_tile_0_2_2),
		.side_3_track_3_out(vertical_tile_1_2_to_tile_0_2_3),
		.side_3_track_0_in(vertical_tile_0_2_to_tile_1_2_0),
		.side_3_track_1_in(vertical_tile_0_2_to_tile_1_2_1),
		.side_3_track_2_in(vertical_tile_0_2_to_tile_1_2_2),
		.side_3_track_3_in(vertical_tile_0_2_to_tile_1_2_3),
		.side_1_track_0_out(vertical_tile_1_2_to_tile_2_2_0),
		.side_1_track_1_out(vertical_tile_1_2_to_tile_2_2_1),
		.side_1_track_2_out(vertical_tile_1_2_to_tile_2_2_2),
		.side_1_track_3_out(vertical_tile_1_2_to_tile_2_2_3),
		.side_1_track_0_in(vertical_tile_2_2_to_tile_1_2_0),
		.side_1_track_1_in(vertical_tile_2_2_to_tile_1_2_1),
		.side_1_track_2_in(vertical_tile_2_2_to_tile_1_2_2),
		.side_1_track_3_in(vertical_tile_2_2_to_tile_1_2_3),
		.side_2_track_0_out(horizontal_tile_1_2_to_tile_1_1_0),
		.side_2_track_1_out(horizontal_tile_1_2_to_tile_1_1_1),
		.side_2_track_2_out(horizontal_tile_1_2_to_tile_1_1_2),
		.side_2_track_3_out(horizontal_tile_1_2_to_tile_1_1_3),
		.side_2_track_0_in(horizontal_tile_1_1_to_tile_1_2_0),
		.side_2_track_1_in(horizontal_tile_1_1_to_tile_1_2_1),
		.side_2_track_2_in(horizontal_tile_1_1_to_tile_1_2_2),
		.side_2_track_3_in(horizontal_tile_1_1_to_tile_1_2_3),
		.side_0_track_0_in(pe_tile_1_2_in_wire_0_0_const),
		.side_0_track_1_in(pe_tile_1_2_in_wire_0_1_const),
		.side_0_track_2_in(pe_tile_1_2_in_wire_0_2_const),
		.side_0_track_3_in(pe_tile_1_2_in_wire_0_3_const),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_1_2_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_0_const_20(
		.out(pe_tile_1_2_in_wire_0_0_const),
		.in(wire_20)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_2_in_wire_0_0_const_20_const(
		.out(wire_20)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_1_const_21(
		.out(pe_tile_1_2_in_wire_0_1_const),
		.in(wire_21)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_2_in_wire_0_1_const_21_const(
		.out(wire_21)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_2_const_22(
		.out(pe_tile_1_2_in_wire_0_2_const),
		.in(wire_22)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_2_in_wire_0_2_const_22_const(
		.out(wire_22)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_3_const_23(
		.out(pe_tile_1_2_in_wire_0_3_const),
		.in(wire_23)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_1_2_in_wire_0_3_const_23_const(
		.out(wire_23)
	);

	assign_mod #(.width(16))  assign_pe_tile_1_2_id_wire_24(
		.out(pe_tile_1_2_id_wire),
		.in(wire_24)
	);

	const_mod #(.value(16'd9), .width(16))  assign_pe_tile_1_2_id_wire_24_const(
		.out(wire_24)
	);

	pe_tile pe_tile_2_0(
		.side_3_track_0_out(vertical_tile_2_0_to_tile_1_0_0),
		.side_3_track_1_out(vertical_tile_2_0_to_tile_1_0_1),
		.side_3_track_2_out(vertical_tile_2_0_to_tile_1_0_2),
		.side_3_track_3_out(vertical_tile_2_0_to_tile_1_0_3),
		.side_3_track_0_in(vertical_tile_1_0_to_tile_2_0_0),
		.side_3_track_1_in(vertical_tile_1_0_to_tile_2_0_1),
		.side_3_track_2_in(vertical_tile_1_0_to_tile_2_0_2),
		.side_3_track_3_in(vertical_tile_1_0_to_tile_2_0_3),
		.side_1_track_0_out(out_pad_0_pin_0_to_pe_tile_2_0_side_1_track_0_out),
		.side_1_track_1_out(out_pad_0_pin_1_to_pe_tile_2_0_side_1_track_1_out),
		.side_1_track_2_out(out_pad_0_pin_2_to_pe_tile_2_0_side_1_track_2_out),
		.side_1_track_3_out(out_pad_0_pin_3_to_pe_tile_2_0_side_1_track_3_out),
		.side_1_track_0_in(pe_tile_2_0_side_1_track_0_in_const),
		.side_1_track_1_in(pe_tile_2_0_side_1_track_1_in_const),
		.side_1_track_2_in(pe_tile_2_0_side_1_track_2_in_const),
		.side_1_track_3_in(pe_tile_2_0_side_1_track_3_in_const),
		.side_2_track_0_in(pe_tile_2_0side_2_track_0_in_const),
		.side_2_track_1_in(pe_tile_2_0side_2_track_1_in_const),
		.side_2_track_2_in(pe_tile_2_0side_2_track_2_in_const),
		.side_2_track_3_in(pe_tile_2_0side_2_track_3_in_const),
		.side_0_track_0_out(horizontal_tile_2_0_to_tile_2_1_0),
		.side_0_track_1_out(horizontal_tile_2_0_to_tile_2_1_1),
		.side_0_track_2_out(horizontal_tile_2_0_to_tile_2_1_2),
		.side_0_track_3_out(horizontal_tile_2_0_to_tile_2_1_3),
		.side_0_track_0_in(horizontal_tile_2_1_to_tile_2_0_0),
		.side_0_track_1_in(horizontal_tile_2_1_to_tile_2_0_1),
		.side_0_track_2_in(horizontal_tile_2_1_to_tile_2_0_2),
		.side_0_track_3_in(horizontal_tile_2_1_to_tile_2_0_3),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_2_0_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_side_1_track_0_in_const_25(
		.out(pe_tile_2_0_side_1_track_0_in_const),
		.in(wire_25)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0_side_1_track_0_in_const_25_const(
		.out(wire_25)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_side_1_track_1_in_const_26(
		.out(pe_tile_2_0_side_1_track_1_in_const),
		.in(wire_26)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0_side_1_track_1_in_const_26_const(
		.out(wire_26)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_side_1_track_2_in_const_27(
		.out(pe_tile_2_0_side_1_track_2_in_const),
		.in(wire_27)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0_side_1_track_2_in_const_27_const(
		.out(wire_27)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_side_1_track_3_in_const_28(
		.out(pe_tile_2_0_side_1_track_3_in_const),
		.in(wire_28)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0_side_1_track_3_in_const_28_const(
		.out(wire_28)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0side_2_track_0_in_const_29(
		.out(pe_tile_2_0side_2_track_0_in_const),
		.in(wire_29)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0side_2_track_0_in_const_29_const(
		.out(wire_29)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0side_2_track_1_in_const_30(
		.out(pe_tile_2_0side_2_track_1_in_const),
		.in(wire_30)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0side_2_track_1_in_const_30_const(
		.out(wire_30)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0side_2_track_2_in_const_31(
		.out(pe_tile_2_0side_2_track_2_in_const),
		.in(wire_31)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0side_2_track_2_in_const_31_const(
		.out(wire_31)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0side_2_track_3_in_const_32(
		.out(pe_tile_2_0side_2_track_3_in_const),
		.in(wire_32)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_0side_2_track_3_in_const_32_const(
		.out(wire_32)
	);

	assign_mod #(.width(16))  assign_pe_tile_2_0_id_wire_33(
		.out(pe_tile_2_0_id_wire),
		.in(wire_33)
	);

	const_mod #(.value(16'd10), .width(16))  assign_pe_tile_2_0_id_wire_33_const(
		.out(wire_33)
	);

	pe_tile pe_tile_2_1(
		.side_3_track_0_out(vertical_tile_2_1_to_tile_1_1_0),
		.side_3_track_1_out(vertical_tile_2_1_to_tile_1_1_1),
		.side_3_track_2_out(vertical_tile_2_1_to_tile_1_1_2),
		.side_3_track_3_out(vertical_tile_2_1_to_tile_1_1_3),
		.side_3_track_0_in(vertical_tile_1_1_to_tile_2_1_0),
		.side_3_track_1_in(vertical_tile_1_1_to_tile_2_1_1),
		.side_3_track_2_in(vertical_tile_1_1_to_tile_2_1_2),
		.side_3_track_3_in(vertical_tile_1_1_to_tile_2_1_3),
		.side_1_track_0_out(out_pad_1_pin_0_to_pe_tile_2_1_side_1_track_0_out),
		.side_1_track_1_out(out_pad_1_pin_1_to_pe_tile_2_1_side_1_track_1_out),
		.side_1_track_2_out(out_pad_1_pin_2_to_pe_tile_2_1_side_1_track_2_out),
		.side_1_track_3_out(out_pad_1_pin_3_to_pe_tile_2_1_side_1_track_3_out),
		.side_1_track_0_in(pe_tile_2_1_side_1_track_0_in_const),
		.side_1_track_1_in(pe_tile_2_1_side_1_track_1_in_const),
		.side_1_track_2_in(pe_tile_2_1_side_1_track_2_in_const),
		.side_1_track_3_in(pe_tile_2_1_side_1_track_3_in_const),
		.side_2_track_0_out(horizontal_tile_2_1_to_tile_2_0_0),
		.side_2_track_1_out(horizontal_tile_2_1_to_tile_2_0_1),
		.side_2_track_2_out(horizontal_tile_2_1_to_tile_2_0_2),
		.side_2_track_3_out(horizontal_tile_2_1_to_tile_2_0_3),
		.side_2_track_0_in(horizontal_tile_2_0_to_tile_2_1_0),
		.side_2_track_1_in(horizontal_tile_2_0_to_tile_2_1_1),
		.side_2_track_2_in(horizontal_tile_2_0_to_tile_2_1_2),
		.side_2_track_3_in(horizontal_tile_2_0_to_tile_2_1_3),
		.side_0_track_0_out(horizontal_tile_2_1_to_tile_2_2_0),
		.side_0_track_1_out(horizontal_tile_2_1_to_tile_2_2_1),
		.side_0_track_2_out(horizontal_tile_2_1_to_tile_2_2_2),
		.side_0_track_3_out(horizontal_tile_2_1_to_tile_2_2_3),
		.side_0_track_0_in(horizontal_tile_2_2_to_tile_2_1_0),
		.side_0_track_1_in(horizontal_tile_2_2_to_tile_2_1_1),
		.side_0_track_2_in(horizontal_tile_2_2_to_tile_2_1_2),
		.side_0_track_3_in(horizontal_tile_2_2_to_tile_2_1_3),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_2_1_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_side_1_track_0_in_const_34(
		.out(pe_tile_2_1_side_1_track_0_in_const),
		.in(wire_34)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_1_side_1_track_0_in_const_34_const(
		.out(wire_34)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_side_1_track_1_in_const_35(
		.out(pe_tile_2_1_side_1_track_1_in_const),
		.in(wire_35)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_1_side_1_track_1_in_const_35_const(
		.out(wire_35)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_side_1_track_2_in_const_36(
		.out(pe_tile_2_1_side_1_track_2_in_const),
		.in(wire_36)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_1_side_1_track_2_in_const_36_const(
		.out(wire_36)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_side_1_track_3_in_const_37(
		.out(pe_tile_2_1_side_1_track_3_in_const),
		.in(wire_37)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_1_side_1_track_3_in_const_37_const(
		.out(wire_37)
	);

	assign_mod #(.width(16))  assign_pe_tile_2_1_id_wire_38(
		.out(pe_tile_2_1_id_wire),
		.in(wire_38)
	);

	const_mod #(.value(16'd11), .width(16))  assign_pe_tile_2_1_id_wire_38_const(
		.out(wire_38)
	);

	pe_tile pe_tile_2_2(
		.side_3_track_0_out(vertical_tile_2_2_to_tile_1_2_0),
		.side_3_track_1_out(vertical_tile_2_2_to_tile_1_2_1),
		.side_3_track_2_out(vertical_tile_2_2_to_tile_1_2_2),
		.side_3_track_3_out(vertical_tile_2_2_to_tile_1_2_3),
		.side_3_track_0_in(vertical_tile_1_2_to_tile_2_2_0),
		.side_3_track_1_in(vertical_tile_1_2_to_tile_2_2_1),
		.side_3_track_2_in(vertical_tile_1_2_to_tile_2_2_2),
		.side_3_track_3_in(vertical_tile_1_2_to_tile_2_2_3),
		.side_1_track_0_out(out_pad_2_pin_0_to_pe_tile_2_2_side_1_track_0_out),
		.side_1_track_1_out(out_pad_2_pin_1_to_pe_tile_2_2_side_1_track_1_out),
		.side_1_track_2_out(out_pad_2_pin_2_to_pe_tile_2_2_side_1_track_2_out),
		.side_1_track_3_out(out_pad_2_pin_3_to_pe_tile_2_2_side_1_track_3_out),
		.side_1_track_0_in(pe_tile_2_2_side_1_track_0_in_const),
		.side_1_track_1_in(pe_tile_2_2_side_1_track_1_in_const),
		.side_1_track_2_in(pe_tile_2_2_side_1_track_2_in_const),
		.side_1_track_3_in(pe_tile_2_2_side_1_track_3_in_const),
		.side_2_track_0_out(horizontal_tile_2_2_to_tile_2_1_0),
		.side_2_track_1_out(horizontal_tile_2_2_to_tile_2_1_1),
		.side_2_track_2_out(horizontal_tile_2_2_to_tile_2_1_2),
		.side_2_track_3_out(horizontal_tile_2_2_to_tile_2_1_3),
		.side_2_track_0_in(horizontal_tile_2_1_to_tile_2_2_0),
		.side_2_track_1_in(horizontal_tile_2_1_to_tile_2_2_1),
		.side_2_track_2_in(horizontal_tile_2_1_to_tile_2_2_2),
		.side_2_track_3_in(horizontal_tile_2_1_to_tile_2_2_3),
		.side_0_track_0_in(pe_tile_2_2_in_wire_0_0_const),
		.side_0_track_1_in(pe_tile_2_2_in_wire_0_1_const),
		.side_0_track_2_in(pe_tile_2_2_in_wire_0_2_const),
		.side_0_track_3_in(pe_tile_2_2_in_wire_0_3_const),
		.clk(clk),
		.rst(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_2_2_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_side_1_track_0_in_const_39(
		.out(pe_tile_2_2_side_1_track_0_in_const),
		.in(wire_39)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_side_1_track_0_in_const_39_const(
		.out(wire_39)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_side_1_track_1_in_const_40(
		.out(pe_tile_2_2_side_1_track_1_in_const),
		.in(wire_40)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_side_1_track_1_in_const_40_const(
		.out(wire_40)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_side_1_track_2_in_const_41(
		.out(pe_tile_2_2_side_1_track_2_in_const),
		.in(wire_41)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_side_1_track_2_in_const_41_const(
		.out(wire_41)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_side_1_track_3_in_const_42(
		.out(pe_tile_2_2_side_1_track_3_in_const),
		.in(wire_42)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_side_1_track_3_in_const_42_const(
		.out(wire_42)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_0_const_43(
		.out(pe_tile_2_2_in_wire_0_0_const),
		.in(wire_43)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_in_wire_0_0_const_43_const(
		.out(wire_43)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_1_const_44(
		.out(pe_tile_2_2_in_wire_0_1_const),
		.in(wire_44)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_in_wire_0_1_const_44_const(
		.out(wire_44)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_2_const_45(
		.out(pe_tile_2_2_in_wire_0_2_const),
		.in(wire_45)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_in_wire_0_2_const_45_const(
		.out(wire_45)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_3_const_46(
		.out(pe_tile_2_2_in_wire_0_3_const),
		.in(wire_46)
	);

	const_mod #(.value(1'b0), .width(1))  assign_pe_tile_2_2_in_wire_0_3_const_46_const(
		.out(wire_46)
	);

	assign_mod #(.width(16))  assign_pe_tile_2_2_id_wire_47(
		.out(pe_tile_2_2_id_wire),
		.in(wire_47)
	);

	const_mod #(.value(16'd12), .width(16))  assign_pe_tile_2_2_id_wire_47_const(
		.out(wire_47)
	);



endmodule